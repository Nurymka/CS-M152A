`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   18:03:37 03/05/2019
// Design Name:   ScoreEvaluation
// Module Name:   /home/ise/XilinxVM/csm152a/whackamole/src/tb/ScoreEvaluation_tb.v
// Project Name:  whackamole
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ScoreEvaluation
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module ScoreEvaluation_tb;

	// Outputs
	//wire ;

	// Instantiate the Unit Under Test (UUT)
	//ScoreEvaluation uut (
	//	.()
	//);

	//initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
	//	#100;
        
		// Add stimulus here

	//end
      
endmodule

